library ieee;
use ieee.std_logic_1164.all;

package MIPS_pkg is

	constant	ROM_ADDR_SIZE	: positive := 6;
	constant	RAM_ADDR_SIZE	: positive := 6;

end package MIPS_pkg;

package body MIPS_pkg is

end package body MIPS_pkg;