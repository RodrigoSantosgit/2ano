library ieee;
use ieee.std_logic_1164.all;

library work;
use work.DisplayUnit_pkg.all;

entity MIPSMultiCycle is
	port(	clk 			: in std_logic;
			reset			: in std_logic;
			cpu_rd		: out std_logic;
			cpu_wr		: out std_logic;
			cpu_addrBus	: out std_logic_vector(31 downto 0);
			cpu_dataBus	: inout std_logic_vector(31 downto 0)
		);
end MIPSMultiCycle;

architecture Struct of MIPSMultiCycle is
-- Signals related to the instruction code
	signal si_instr : std_logic_vector(31 downto 0);
	signal si_opcode, si_funct : std_logic_vector(5 downto 0);
	signal si_rs, si_rt, si_rd, si_writeReg : std_logic_vector(4 downto 0);
	signal si_imm : std_logic_vector(15 downto 0);
	signal si_jAddr : std_logic_vector(25 downto 0);
	signal si_offset32, si_left2 : std_logic_vector(31 downto 0);
	
-- Other signals
	signal s_zero : std_logic;
	signal s_pc : std_logic_vector(31 downto 0);
	signal s_aluOper : std_logic_vector(2 downto 0);

-- Data signals
	signal sd_readData1, sd_readData2 : std_logic_vector(31 downto 0);
	signal sd_regA, sd_regB : std_logic_vector(31 downto 0);
	signal sd_aluA, sd_aluB : std_logic_vector(31 downto 0);
	signal sd_aluRes : std_logic_vector(31 downto 0);
	signal sd_aluOut : std_logic_vector(31 downto 0);
	signal sd_data : std_logic_vector(31 downto 0);
	signal sd_writeData : std_logic_vector(31 downto 0);
	
-- Control signals (generated by the control unit)
	signal sc_IorD, sc_RegDst, sc_MemToReg : std_logic;
	signal sc_AluSel_a : std_logic;
	signal sc_AluSel_b, sc_AluOp : std_logic_vector(1 downto 0);	
	signal sc_RegWrite, sc_IrWrite  : std_logic;
	signal sc_PCWrite, sc_PCWriteCond : std_logic;
	signal sc_PCSource : std_logic_vector(1 downto 0);	
	
begin

-- PC update
pcupd:	entity work.PCupdate(Behavioral)	
			port map(clk			=> s_clk,
						reset			=> s_reset,
						zero			=> s_zero,
						PCSource		=> sc_PCSource, 
						PCWrite		=> sc_PCWrite,
						PCWriteCond	=> sc_PCWriteCond,
						PC4			=> sd_aluOut,
						BTA			=> sd_,
						jAddr			=> si_jAddr,
						pc				=> s_pc);

-- MUX M1 (address multiplexer)
mux_m1:	entity work.MUX21_N(Behavioral)
			generic map(N => )
			port map(In0	=> ,
						In1	=> ,
						Sel	=> ,
						MuxOut=> cpu_addrBus);	-- CPU Address Bus		
					
-- Instruction Register
instReg:	entity work.Register_N(Behavioral)
			port map(clk		=> ,
						enable	=> ,
						valIn		=> cpu_dataBus,
						valOut	=> );

-- Data Register
dataReg:	entity work.Register_N(Behavioral)
			port map(clk		=> ,
						enable	=> '1',
						valIn		=> cpu_dataBus,	-- CPU Data Bus
						valOut	=> );
						
-- Splitter
spliter:	entity work.InstSplitter(Behavioral)
			port map(instruction	=> ,
						opcode		=> ,
						rs				=> ,
						rt				=> ,
						rd				=> ,
						funct			=> ,
						imm			=> ,
						jAddr			=> );

-- MUX M2 (Destination register multiplexer)
mux_m2:	entity work.MUX21_N(Behavioral)
			generic map(N => )
			port map(In0	=> ,
						In1	=> ,
						Sel	=> ,
						MuxOut=> );		

-- MUX M3 (Register write data multiplexer)
mux_m3:	entity work.MUX21_N(Behavioral)
			generic map(N => )
			port map(In0	=> ,
						In1	=> ,
						Sel	=> ,
						MuxOut=> );		
						
-- Register File
regfile:	entity work.RegFile(Structural)
			port map(clk			=> clk,
						writeEnable	=> ,
						writeReg		=> ,
						writeData	=> ,
						readReg1		=> ,
						readReg2		=> ,
						readData1	=> ,
						readData2	=> );

-- A Register
regA:	entity work.Register_N(Behavioral)
			port map(clk		=> ,
						enable	=> '1',
						valIn		=> ,
						valOut	=> );

-- B Register
regB:	entity work.Register_N(Behavioral)
			port map(clk		=> ,
						enable	=> '1',
						valIn		=> ,
						valOut	=> );

-- MUX M4 (ALU operand A multiplexer)
mux_m4:	entity work.MUX21_N(Behavioral)
			generic map(N => )
			port map(In0	=> ,
						In1	=> ,
						Sel	=> ,
						MuxOut=> );

-- MUX M5 (ALU operand B multiplexer)
mux_m5:	entity work.MUX41_N(Behavioral)
			generic map(N => )
			port map(In0	=> ,
						In1	=> ,
						In2 	=> ,
						In3 	=> ,
						Sel	=> ,
						MuxOut=> );
						
-- ALU
alu:		entity work.alu32(Behavioral)
			port map(a		=> ,
						b  	=> ,
						oper	=> ,
						res	=> ,
						zero	=> );
						
-- ALU Control		
alucntl:	entity work.ALUControlUnit(Behavioral)
			port map(ALUop		 => ,
						funct		 => ,
						ALUcontrol=> );
						
-- ALUOut Register
regALU:	entity work.Register_N(Behavioral)
			port map(clk		=> ,
						enable	=> '1',
						valIn		=> ,
						valOut	=> );
												
-- left shifter
ls2:		entity work.LeftShifter2(Behavioral)
			port map(dataIn	=> ,
						dataOut	=> );
						
-- sign extend
signext:	entity work.SignExtend(Behavioral)
			port map(dataIn	=> ,
						dataOut	=> );
						
-- Control Unit											
control:	entity work.ControlUnit(Behavioral)
			port map(Clk			=> ,
						Reset			=> ,
						OpCode 		=> ,
						PCWrite		=> sc_PCWrite,
						IRWrite		=> sc_IrWrite,
						IorD			=> sc_IorD,
						PCSource		=> sc_PCSource,
						RegDest		=> sc_RegDst,
						PCWriteCond	=> sc_PCWriteCond,
						MemRead		=> cpu_rd,			-- CPU read signal
						MemWrite		=> cpu_wr,			-- CPU write signal
						MemToReg		=> sc_MemToReg,
						ALUSelA		=> sc_AluSel_a,
						ALUSelB		=> sc_AluSel_b,
						RegWrite		=> sc_RegWrite,
						ALUop 		=> sc_AluOp);

-- Tri-state logic (data bus)
	cpu_dataBus <= sd_regB when cpu_wr = '1' else (others => 'Z');	-- CPU cpu_dataBus
	
-- Connection to DisplayUnit (ALU result, shown as Instr. Memory Data)
	DU_IMdata <= sd_aluRes;
						
end Struct;

